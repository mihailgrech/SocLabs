module vl1(x);
output x;

assign x = 1'b1;
endmodule
