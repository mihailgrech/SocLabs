module vl2(y);
output y;

assign y = 1'b0;
endmodule
