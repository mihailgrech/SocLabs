module decoder(Q, AG);
  input [3:0] Q;
  output [6:0] AG;
  reg [6:0] AG;
  
  always @(Q)
    case (Q)
      4'b0000: AG = 7'b1111110;
      4'b0001: AG = 7'b0110000;
      4'b0010: AG = 7'b1101101;
      4'b0011: AG = 7'b1111001;
      4'b0100: AG = 7'b0110011;
      4'b0101: AG = 7'b1011011;
      4'b0110: AG = 7'b1011111;
      4'b0111: AG = 7'b1110000;
      4'b1000: AG = 7'b1111111;
      4'b1001: AG = 7'b1111011;
      4'b1010: AG = 7'b1110111;
      4'b1011: AG = 7'b0011111;
      4'b1100: AG = 7'b1001110;
      4'b1101: AG = 7'b0111101;
      4'b1110: AG = 7'b1001111;
      4'b1111: AG = 7'b1000111;
    endcase
    
endmodule